LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY ROM IS
	PORT(
		entrada : IN  STD_LOGIC_VECTOR (7 DOWNTO 0);
		saida	: OUT STD_LOGIC_VECTOR (7 DOWNTO 0));
END ROM;

ARCHITECTURE arch OF ROM IS
BEGIN
	WITH entrada SELECT
	--  saida <=    "DADO_MEM" WHEN "ADDR_MEM",
		saida <= 	"00101111" WHEN "00000000",	-- LDA
					"00000000" WHEN "00000001", -- 0x00
					"01010000" WHEN "00000010", -- AND
					"00001111" WHEN "00000011", -- 0x0F
					"00000000" WHEN "00000100", -- NOP
					"10000000" WHEN "00000101", -- JMP
					"00000000" WHEN "00000110", -- 0x00
					"00000000" WHEN OTHERS;
END arch; 